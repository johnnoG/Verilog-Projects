`include "and.sv"
`include "nor.sv"
`include "xor.sv"
`include "mux.sv"
`include "fas.sv"
`include "alu.sv"