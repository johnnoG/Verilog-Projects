// Code your testbench here
// or browse Examples

`include "demo.sv"
`include "mux4_tb.sv"
`include "rip_fas_tb.sv"
`include "alu_4bit_tb_sv"
